library verilog;
use verilog.vl_types.all;
entity cyclone_pll is
    generic(
        operation_mode  : string  := "normal";
        qualify_conf_done: string  := "off";
        compensate_clock: string  := "clk0";
        pll_type        : string  := "auto";
        scan_chain      : string  := "long";
        lpm_type        : string  := "cyclone_pll";
        clk0_multiply_by: integer := 1;
        clk0_divide_by  : integer := 1;
        clk0_phase_shift: integer := 0;
        clk0_time_delay : integer := 0;
        clk0_duty_cycle : integer := 50;
        clk1_multiply_by: integer := 1;
        clk1_divide_by  : integer := 1;
        clk1_phase_shift: integer := 0;
        clk1_time_delay : integer := 0;
        clk1_duty_cycle : integer := 50;
        clk2_multiply_by: integer := 1;
        clk2_divide_by  : integer := 1;
        clk2_phase_shift: integer := 0;
        clk2_time_delay : integer := 0;
        clk2_duty_cycle : integer := 50;
        clk3_multiply_by: integer := 1;
        clk3_divide_by  : integer := 1;
        clk3_phase_shift: integer := 0;
        clk3_time_delay : integer := 0;
        clk3_duty_cycle : integer := 50;
        clk4_multiply_by: integer := 1;
        clk4_divide_by  : integer := 1;
        clk4_phase_shift: integer := 0;
        clk4_time_delay : integer := 0;
        clk4_duty_cycle : integer := 50;
        clk5_multiply_by: integer := 1;
        clk5_divide_by  : integer := 1;
        clk5_phase_shift: integer := 0;
        clk5_time_delay : integer := 0;
        clk5_duty_cycle : integer := 50;
        extclk0_multiply_by: integer := 1;
        extclk0_divide_by: integer := 1;
        extclk0_phase_shift: integer := 0;
        extclk0_time_delay: integer := 0;
        extclk0_duty_cycle: integer := 50;
        extclk1_multiply_by: integer := 1;
        extclk1_divide_by: integer := 1;
        extclk1_phase_shift: integer := 0;
        extclk1_time_delay: integer := 0;
        extclk1_duty_cycle: integer := 50;
        extclk2_multiply_by: integer := 1;
        extclk2_divide_by: integer := 1;
        extclk2_phase_shift: integer := 0;
        extclk2_time_delay: integer := 0;
        extclk2_duty_cycle: integer := 50;
        extclk3_multiply_by: integer := 1;
        extclk3_divide_by: integer := 1;
        extclk3_phase_shift: integer := 0;
        extclk3_time_delay: integer := 0;
        extclk3_duty_cycle: integer := 50;
        primary_clock   : string  := "inclk0";
        inclk0_input_frequency: integer := 10000;
        inclk1_input_frequency: integer := 10000;
        gate_lock_signal: string  := "no";
        gate_lock_counter: integer := 1;
        valid_lock_multiplier: integer := 5;
        invalid_lock_multiplier: integer := 5;
        switch_over_on_lossclk: string  := "off";
        switch_over_on_gated_lock: string  := "off";
        switch_over_counter: integer := 1;
        enable_switch_over_counter: string  := "off";
        feedback_source : string  := "extclk0";
        bandwidth       : integer := 0;
        bandwidth_type  : string  := "auto";
        spread_frequency: integer := 0;
        common_rx_tx    : string  := "off";
        rx_outclock_resource: string  := "auto";
        use_vco_bypass  : string  := "false";
        use_dc_coupling : string  := "false";
        pfd_min         : integer := 0;
        pfd_max         : integer := 0;
        vco_min         : integer := 0;
        vco_max         : integer := 0;
        vco_center      : integer := 0;
        m_initial       : integer := 1;
        m               : integer := 0;
        n               : integer := 1;
        m2              : integer := 1;
        n2              : integer := 1;
        ss              : integer := 0;
        l0_high         : integer := 1;
        l0_low          : integer := 1;
        l0_initial      : integer := 1;
        l0_mode         : string  := "bypass";
        l0_ph           : integer := 0;
        l0_time_delay   : integer := 0;
        l1_high         : integer := 1;
        l1_low          : integer := 1;
        l1_initial      : integer := 1;
        l1_mode         : string  := "bypass";
        l1_ph           : integer := 0;
        l1_time_delay   : integer := 0;
        g0_high         : integer := 1;
        g0_low          : integer := 1;
        g0_initial      : integer := 1;
        g0_mode         : string  := "bypass";
        g0_ph           : integer := 0;
        g0_time_delay   : integer := 0;
        g1_high         : integer := 1;
        g1_low          : integer := 1;
        g1_initial      : integer := 1;
        g1_mode         : string  := "bypass";
        g1_ph           : integer := 0;
        g1_time_delay   : integer := 0;
        g2_high         : integer := 1;
        g2_low          : integer := 1;
        g2_initial      : integer := 1;
        g2_mode         : string  := "bypass";
        g2_ph           : integer := 0;
        g2_time_delay   : integer := 0;
        g3_high         : integer := 1;
        g3_low          : integer := 1;
        g3_initial      : integer := 1;
        g3_mode         : string  := "bypass";
        g3_ph           : integer := 0;
        g3_time_delay   : integer := 0;
        e0_high         : integer := 1;
        e0_low          : integer := 1;
        e0_initial      : integer := 1;
        e0_mode         : string  := "bypass";
        e0_ph           : integer := 0;
        e0_time_delay   : integer := 0;
        e1_high         : integer := 1;
        e1_low          : integer := 1;
        e1_initial      : integer := 1;
        e1_mode         : string  := "bypass";
        e1_ph           : integer := 0;
        e1_time_delay   : integer := 0;
        e2_high         : integer := 1;
        e2_low          : integer := 1;
        e2_initial      : integer := 1;
        e2_mode         : string  := "bypass";
        e2_ph           : integer := 0;
        e2_time_delay   : integer := 0;
        e3_high         : integer := 1;
        e3_low          : integer := 1;
        e3_initial      : integer := 1;
        e3_mode         : string  := "bypass";
        e3_ph           : integer := 0;
        e3_time_delay   : integer := 0;
        m_ph            : integer := 0;
        m_time_delay    : integer := 0;
        n_time_delay    : integer := 0;
        extclk0_counter : string  := "e0";
        extclk1_counter : string  := "e1";
        extclk2_counter : string  := "e2";
        extclk3_counter : string  := "e3";
        clk0_counter    : string  := "g0";
        clk1_counter    : string  := "g1";
        clk2_counter    : string  := "g2";
        clk3_counter    : string  := "g3";
        clk4_counter    : string  := "l0";
        clk5_counter    : string  := "l1";
        enable0_counter : string  := "l0";
        enable1_counter : string  := "l0";
        charge_pump_current: integer := 0;
        loop_filter_r   : string  := "1.0";
        loop_filter_c   : integer := 1;
        pll_compensation_delay: integer := 0;
        simulation_type : string  := "timing";
        source_is_pll   : string  := "off";
        down_spread     : string  := "0.0";
        clk0_phase_shift_num: integer := 0;
        clk1_phase_shift_num: integer := 0;
        clk2_phase_shift_num: integer := 0;
        family_name     : string  := "Cyclone";
        skip_vco        : string  := "off";
        clk0_use_even_counter_mode: string  := "off";
        clk1_use_even_counter_mode: string  := "off";
        clk2_use_even_counter_mode: string  := "off";
        clk3_use_even_counter_mode: string  := "off";
        clk4_use_even_counter_mode: string  := "off";
        clk5_use_even_counter_mode: string  := "off";
        extclk0_use_even_counter_mode: string  := "off";
        extclk1_use_even_counter_mode: string  := "off";
        extclk2_use_even_counter_mode: string  := "off";
        extclk3_use_even_counter_mode: string  := "off";
        clk0_use_even_counter_value: string  := "off";
        clk1_use_even_counter_value: string  := "off";
        clk2_use_even_counter_value: string  := "off";
        clk3_use_even_counter_value: string  := "off";
        clk4_use_even_counter_value: string  := "off";
        clk5_use_even_counter_value: string  := "off";
        extclk0_use_even_counter_value: string  := "off";
        extclk1_use_even_counter_value: string  := "off";
        extclk2_use_even_counter_value: string  := "off";
        extclk3_use_even_counter_value: string  := "off";
        EGPP_SCAN_CHAIN : integer := 289;
        GPP_SCAN_CHAIN  : integer := 193;
        TRST            : integer := 5000;
        TRSTCLK         : integer := 5000
    );
    port(
        inclk           : in     vl_logic_vector(1 downto 0);
        fbin            : in     vl_logic;
        ena             : in     vl_logic;
        clkswitch       : in     vl_logic;
        areset          : in     vl_logic;
        pfdena          : in     vl_logic;
        clkena          : in     vl_logic_vector(5 downto 0);
        extclkena       : in     vl_logic_vector(3 downto 0);
        scanclk         : in     vl_logic;
        scanaclr        : in     vl_logic;
        scandata        : in     vl_logic;
        clk             : out    vl_logic_vector(5 downto 0);
        extclk          : out    vl_logic_vector(3 downto 0);
        clkbad          : out    vl_logic_vector(1 downto 0);
        activeclock     : out    vl_logic;
        locked          : out    vl_logic;
        clkloss         : out    vl_logic;
        scandataout     : out    vl_logic;
        comparator      : in     vl_logic;
        enable0         : out    vl_logic;
        enable1         : out    vl_logic
    );
    attribute mti_svvh_generic_type : integer;
    attribute mti_svvh_generic_type of operation_mode : constant is 1;
    attribute mti_svvh_generic_type of qualify_conf_done : constant is 1;
    attribute mti_svvh_generic_type of compensate_clock : constant is 1;
    attribute mti_svvh_generic_type of pll_type : constant is 1;
    attribute mti_svvh_generic_type of scan_chain : constant is 1;
    attribute mti_svvh_generic_type of lpm_type : constant is 1;
    attribute mti_svvh_generic_type of clk0_multiply_by : constant is 1;
    attribute mti_svvh_generic_type of clk0_divide_by : constant is 1;
    attribute mti_svvh_generic_type of clk0_phase_shift : constant is 1;
    attribute mti_svvh_generic_type of clk0_time_delay : constant is 1;
    attribute mti_svvh_generic_type of clk0_duty_cycle : constant is 1;
    attribute mti_svvh_generic_type of clk1_multiply_by : constant is 1;
    attribute mti_svvh_generic_type of clk1_divide_by : constant is 1;
    attribute mti_svvh_generic_type of clk1_phase_shift : constant is 1;
    attribute mti_svvh_generic_type of clk1_time_delay : constant is 1;
    attribute mti_svvh_generic_type of clk1_duty_cycle : constant is 1;
    attribute mti_svvh_generic_type of clk2_multiply_by : constant is 1;
    attribute mti_svvh_generic_type of clk2_divide_by : constant is 1;
    attribute mti_svvh_generic_type of clk2_phase_shift : constant is 1;
    attribute mti_svvh_generic_type of clk2_time_delay : constant is 1;
    attribute mti_svvh_generic_type of clk2_duty_cycle : constant is 1;
    attribute mti_svvh_generic_type of clk3_multiply_by : constant is 1;
    attribute mti_svvh_generic_type of clk3_divide_by : constant is 1;
    attribute mti_svvh_generic_type of clk3_phase_shift : constant is 1;
    attribute mti_svvh_generic_type of clk3_time_delay : constant is 1;
    attribute mti_svvh_generic_type of clk3_duty_cycle : constant is 1;
    attribute mti_svvh_generic_type of clk4_multiply_by : constant is 1;
    attribute mti_svvh_generic_type of clk4_divide_by : constant is 1;
    attribute mti_svvh_generic_type of clk4_phase_shift : constant is 1;
    attribute mti_svvh_generic_type of clk4_time_delay : constant is 1;
    attribute mti_svvh_generic_type of clk4_duty_cycle : constant is 1;
    attribute mti_svvh_generic_type of clk5_multiply_by : constant is 1;
    attribute mti_svvh_generic_type of clk5_divide_by : constant is 1;
    attribute mti_svvh_generic_type of clk5_phase_shift : constant is 1;
    attribute mti_svvh_generic_type of clk5_time_delay : constant is 1;
    attribute mti_svvh_generic_type of clk5_duty_cycle : constant is 1;
    attribute mti_svvh_generic_type of extclk0_multiply_by : constant is 1;
    attribute mti_svvh_generic_type of extclk0_divide_by : constant is 1;
    attribute mti_svvh_generic_type of extclk0_phase_shift : constant is 1;
    attribute mti_svvh_generic_type of extclk0_time_delay : constant is 1;
    attribute mti_svvh_generic_type of extclk0_duty_cycle : constant is 1;
    attribute mti_svvh_generic_type of extclk1_multiply_by : constant is 1;
    attribute mti_svvh_generic_type of extclk1_divide_by : constant is 1;
    attribute mti_svvh_generic_type of extclk1_phase_shift : constant is 1;
    attribute mti_svvh_generic_type of extclk1_time_delay : constant is 1;
    attribute mti_svvh_generic_type of extclk1_duty_cycle : constant is 1;
    attribute mti_svvh_generic_type of extclk2_multiply_by : constant is 1;
    attribute mti_svvh_generic_type of extclk2_divide_by : constant is 1;
    attribute mti_svvh_generic_type of extclk2_phase_shift : constant is 1;
    attribute mti_svvh_generic_type of extclk2_time_delay : constant is 1;
    attribute mti_svvh_generic_type of extclk2_duty_cycle : constant is 1;
    attribute mti_svvh_generic_type of extclk3_multiply_by : constant is 1;
    attribute mti_svvh_generic_type of extclk3_divide_by : constant is 1;
    attribute mti_svvh_generic_type of extclk3_phase_shift : constant is 1;
    attribute mti_svvh_generic_type of extclk3_time_delay : constant is 1;
    attribute mti_svvh_generic_type of extclk3_duty_cycle : constant is 1;
    attribute mti_svvh_generic_type of primary_clock : constant is 1;
    attribute mti_svvh_generic_type of inclk0_input_frequency : constant is 1;
    attribute mti_svvh_generic_type of inclk1_input_frequency : constant is 1;
    attribute mti_svvh_generic_type of gate_lock_signal : constant is 1;
    attribute mti_svvh_generic_type of gate_lock_counter : constant is 1;
    attribute mti_svvh_generic_type of valid_lock_multiplier : constant is 1;
    attribute mti_svvh_generic_type of invalid_lock_multiplier : constant is 1;
    attribute mti_svvh_generic_type of switch_over_on_lossclk : constant is 1;
    attribute mti_svvh_generic_type of switch_over_on_gated_lock : constant is 1;
    attribute mti_svvh_generic_type of switch_over_counter : constant is 1;
    attribute mti_svvh_generic_type of enable_switch_over_counter : constant is 1;
    attribute mti_svvh_generic_type of feedback_source : constant is 1;
    attribute mti_svvh_generic_type of bandwidth : constant is 1;
    attribute mti_svvh_generic_type of bandwidth_type : constant is 1;
    attribute mti_svvh_generic_type of spread_frequency : constant is 1;
    attribute mti_svvh_generic_type of common_rx_tx : constant is 1;
    attribute mti_svvh_generic_type of rx_outclock_resource : constant is 1;
    attribute mti_svvh_generic_type of use_vco_bypass : constant is 1;
    attribute mti_svvh_generic_type of use_dc_coupling : constant is 1;
    attribute mti_svvh_generic_type of pfd_min : constant is 1;
    attribute mti_svvh_generic_type of pfd_max : constant is 1;
    attribute mti_svvh_generic_type of vco_min : constant is 1;
    attribute mti_svvh_generic_type of vco_max : constant is 1;
    attribute mti_svvh_generic_type of vco_center : constant is 1;
    attribute mti_svvh_generic_type of m_initial : constant is 1;
    attribute mti_svvh_generic_type of m : constant is 1;
    attribute mti_svvh_generic_type of n : constant is 1;
    attribute mti_svvh_generic_type of m2 : constant is 1;
    attribute mti_svvh_generic_type of n2 : constant is 1;
    attribute mti_svvh_generic_type of ss : constant is 1;
    attribute mti_svvh_generic_type of l0_high : constant is 1;
    attribute mti_svvh_generic_type of l0_low : constant is 1;
    attribute mti_svvh_generic_type of l0_initial : constant is 1;
    attribute mti_svvh_generic_type of l0_mode : constant is 1;
    attribute mti_svvh_generic_type of l0_ph : constant is 1;
    attribute mti_svvh_generic_type of l0_time_delay : constant is 1;
    attribute mti_svvh_generic_type of l1_high : constant is 1;
    attribute mti_svvh_generic_type of l1_low : constant is 1;
    attribute mti_svvh_generic_type of l1_initial : constant is 1;
    attribute mti_svvh_generic_type of l1_mode : constant is 1;
    attribute mti_svvh_generic_type of l1_ph : constant is 1;
    attribute mti_svvh_generic_type of l1_time_delay : constant is 1;
    attribute mti_svvh_generic_type of g0_high : constant is 1;
    attribute mti_svvh_generic_type of g0_low : constant is 1;
    attribute mti_svvh_generic_type of g0_initial : constant is 1;
    attribute mti_svvh_generic_type of g0_mode : constant is 1;
    attribute mti_svvh_generic_type of g0_ph : constant is 1;
    attribute mti_svvh_generic_type of g0_time_delay : constant is 1;
    attribute mti_svvh_generic_type of g1_high : constant is 1;
    attribute mti_svvh_generic_type of g1_low : constant is 1;
    attribute mti_svvh_generic_type of g1_initial : constant is 1;
    attribute mti_svvh_generic_type of g1_mode : constant is 1;
    attribute mti_svvh_generic_type of g1_ph : constant is 1;
    attribute mti_svvh_generic_type of g1_time_delay : constant is 1;
    attribute mti_svvh_generic_type of g2_high : constant is 1;
    attribute mti_svvh_generic_type of g2_low : constant is 1;
    attribute mti_svvh_generic_type of g2_initial : constant is 1;
    attribute mti_svvh_generic_type of g2_mode : constant is 1;
    attribute mti_svvh_generic_type of g2_ph : constant is 1;
    attribute mti_svvh_generic_type of g2_time_delay : constant is 1;
    attribute mti_svvh_generic_type of g3_high : constant is 1;
    attribute mti_svvh_generic_type of g3_low : constant is 1;
    attribute mti_svvh_generic_type of g3_initial : constant is 1;
    attribute mti_svvh_generic_type of g3_mode : constant is 1;
    attribute mti_svvh_generic_type of g3_ph : constant is 1;
    attribute mti_svvh_generic_type of g3_time_delay : constant is 1;
    attribute mti_svvh_generic_type of e0_high : constant is 1;
    attribute mti_svvh_generic_type of e0_low : constant is 1;
    attribute mti_svvh_generic_type of e0_initial : constant is 1;
    attribute mti_svvh_generic_type of e0_mode : constant is 1;
    attribute mti_svvh_generic_type of e0_ph : constant is 1;
    attribute mti_svvh_generic_type of e0_time_delay : constant is 1;
    attribute mti_svvh_generic_type of e1_high : constant is 1;
    attribute mti_svvh_generic_type of e1_low : constant is 1;
    attribute mti_svvh_generic_type of e1_initial : constant is 1;
    attribute mti_svvh_generic_type of e1_mode : constant is 1;
    attribute mti_svvh_generic_type of e1_ph : constant is 1;
    attribute mti_svvh_generic_type of e1_time_delay : constant is 1;
    attribute mti_svvh_generic_type of e2_high : constant is 1;
    attribute mti_svvh_generic_type of e2_low : constant is 1;
    attribute mti_svvh_generic_type of e2_initial : constant is 1;
    attribute mti_svvh_generic_type of e2_mode : constant is 1;
    attribute mti_svvh_generic_type of e2_ph : constant is 1;
    attribute mti_svvh_generic_type of e2_time_delay : constant is 1;
    attribute mti_svvh_generic_type of e3_high : constant is 1;
    attribute mti_svvh_generic_type of e3_low : constant is 1;
    attribute mti_svvh_generic_type of e3_initial : constant is 1;
    attribute mti_svvh_generic_type of e3_mode : constant is 1;
    attribute mti_svvh_generic_type of e3_ph : constant is 1;
    attribute mti_svvh_generic_type of e3_time_delay : constant is 1;
    attribute mti_svvh_generic_type of m_ph : constant is 1;
    attribute mti_svvh_generic_type of m_time_delay : constant is 1;
    attribute mti_svvh_generic_type of n_time_delay : constant is 1;
    attribute mti_svvh_generic_type of extclk0_counter : constant is 1;
    attribute mti_svvh_generic_type of extclk1_counter : constant is 1;
    attribute mti_svvh_generic_type of extclk2_counter : constant is 1;
    attribute mti_svvh_generic_type of extclk3_counter : constant is 1;
    attribute mti_svvh_generic_type of clk0_counter : constant is 1;
    attribute mti_svvh_generic_type of clk1_counter : constant is 1;
    attribute mti_svvh_generic_type of clk2_counter : constant is 1;
    attribute mti_svvh_generic_type of clk3_counter : constant is 1;
    attribute mti_svvh_generic_type of clk4_counter : constant is 1;
    attribute mti_svvh_generic_type of clk5_counter : constant is 1;
    attribute mti_svvh_generic_type of enable0_counter : constant is 1;
    attribute mti_svvh_generic_type of enable1_counter : constant is 1;
    attribute mti_svvh_generic_type of charge_pump_current : constant is 1;
    attribute mti_svvh_generic_type of loop_filter_r : constant is 1;
    attribute mti_svvh_generic_type of loop_filter_c : constant is 1;
    attribute mti_svvh_generic_type of pll_compensation_delay : constant is 1;
    attribute mti_svvh_generic_type of simulation_type : constant is 1;
    attribute mti_svvh_generic_type of source_is_pll : constant is 1;
    attribute mti_svvh_generic_type of down_spread : constant is 1;
    attribute mti_svvh_generic_type of clk0_phase_shift_num : constant is 1;
    attribute mti_svvh_generic_type of clk1_phase_shift_num : constant is 1;
    attribute mti_svvh_generic_type of clk2_phase_shift_num : constant is 1;
    attribute mti_svvh_generic_type of family_name : constant is 1;
    attribute mti_svvh_generic_type of skip_vco : constant is 1;
    attribute mti_svvh_generic_type of clk0_use_even_counter_mode : constant is 1;
    attribute mti_svvh_generic_type of clk1_use_even_counter_mode : constant is 1;
    attribute mti_svvh_generic_type of clk2_use_even_counter_mode : constant is 1;
    attribute mti_svvh_generic_type of clk3_use_even_counter_mode : constant is 1;
    attribute mti_svvh_generic_type of clk4_use_even_counter_mode : constant is 1;
    attribute mti_svvh_generic_type of clk5_use_even_counter_mode : constant is 1;
    attribute mti_svvh_generic_type of extclk0_use_even_counter_mode : constant is 1;
    attribute mti_svvh_generic_type of extclk1_use_even_counter_mode : constant is 1;
    attribute mti_svvh_generic_type of extclk2_use_even_counter_mode : constant is 1;
    attribute mti_svvh_generic_type of extclk3_use_even_counter_mode : constant is 1;
    attribute mti_svvh_generic_type of clk0_use_even_counter_value : constant is 1;
    attribute mti_svvh_generic_type of clk1_use_even_counter_value : constant is 1;
    attribute mti_svvh_generic_type of clk2_use_even_counter_value : constant is 1;
    attribute mti_svvh_generic_type of clk3_use_even_counter_value : constant is 1;
    attribute mti_svvh_generic_type of clk4_use_even_counter_value : constant is 1;
    attribute mti_svvh_generic_type of clk5_use_even_counter_value : constant is 1;
    attribute mti_svvh_generic_type of extclk0_use_even_counter_value : constant is 1;
    attribute mti_svvh_generic_type of extclk1_use_even_counter_value : constant is 1;
    attribute mti_svvh_generic_type of extclk2_use_even_counter_value : constant is 1;
    attribute mti_svvh_generic_type of extclk3_use_even_counter_value : constant is 1;
    attribute mti_svvh_generic_type of EGPP_SCAN_CHAIN : constant is 1;
    attribute mti_svvh_generic_type of GPP_SCAN_CHAIN : constant is 1;
    attribute mti_svvh_generic_type of TRST : constant is 1;
    attribute mti_svvh_generic_type of TRSTCLK : constant is 1;
end cyclone_pll;

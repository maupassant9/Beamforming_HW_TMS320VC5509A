library verilog;
use verilog.vl_types.all;
entity altsyncram is
    generic(
        width_a         : integer := 1;
        widthad_a       : integer := 1;
        numwords_a      : integer := 0;
        outdata_reg_a   : string  := "UNREGISTERED";
        address_aclr_a  : string  := "NONE";
        outdata_aclr_a  : string  := "NONE";
        indata_aclr_a   : string  := "NONE";
        wrcontrol_aclr_a: string  := "NONE";
        byteena_aclr_a  : string  := "NONE";
        width_byteena_a : integer := 1;
        width_b         : integer := 1;
        widthad_b       : integer := 1;
        numwords_b      : integer := 0;
        rdcontrol_reg_b : string  := "CLOCK1";
        address_reg_b   : string  := "CLOCK1";
        outdata_reg_b   : string  := "UNREGISTERED";
        outdata_aclr_b  : string  := "NONE";
        rdcontrol_aclr_b: string  := "NONE";
        indata_reg_b    : string  := "CLOCK1";
        wrcontrol_wraddress_reg_b: string  := "CLOCK1";
        byteena_reg_b   : string  := "CLOCK1";
        indata_aclr_b   : string  := "NONE";
        wrcontrol_aclr_b: string  := "NONE";
        address_aclr_b  : string  := "NONE";
        byteena_aclr_b  : string  := "NONE";
        width_byteena_b : integer := 1;
        clock_enable_input_a: string  := "NORMAL";
        clock_enable_output_a: string  := "NORMAL";
        clock_enable_input_b: string  := "NORMAL";
        clock_enable_output_b: string  := "NORMAL";
        clock_enable_core_a: string  := "USE_INPUT_CLKEN";
        clock_enable_core_b: string  := "USE_INPUT_CLKEN";
        read_during_write_mode_port_a: string  := "NEW_DATA_NO_NBE_READ";
        read_during_write_mode_port_b: string  := "NEW_DATA_NO_NBE_READ";
        enable_ecc      : string  := "FALSE";
        width_eccstatus : integer := 3;
        ecc_pipeline_stage_enabled: string  := "FALSE";
        operation_mode  : string  := "BIDIR_DUAL_PORT";
        byte_size       : integer := 0;
        read_during_write_mode_mixed_ports: string  := "DONT_CARE";
        ram_block_type  : string  := "AUTO";
        init_file       : string  := "UNUSED";
        init_file_layout: string  := "UNUSED";
        maximum_depth   : integer := 0;
        intended_device_family: string  := "Stratix";
        lpm_hint        : string  := "UNUSED";
        lpm_type        : string  := "altsyncram";
        implement_in_les: string  := "OFF";
        power_up_uninitialized: string  := "FALSE";
        sim_show_memory_data_in_port_b_layout: string  := "OFF";
        is_lutram       : vl_notype;
        is_bidir_and_wrcontrol_addb_clk0: vl_notype;
        is_bidir_and_wrcontrol_addb_clk1: vl_notype;
        check_simultaneous_read_write: vl_notype;
        dual_port_addreg_b_clk0: vl_notype;
        dual_port_addreg_b_clk1: vl_notype;
        i_byte_size_tmp : vl_notype;
        i_lutram_read   : vl_notype;
        enable_mem_data_b_reading: vl_notype;
        family_arriav   : vl_notype;
        family_cyclonev : vl_notype;
        family_base_arriav: vl_notype;
        family_stratixvi: vl_notype;
        family_arriavi  : vl_notype;
        family_nightfury: vl_notype;
        family_arriavgz : vl_notype;
        family_stratixv : vl_notype;
        family_hardcopyiv: vl_notype;
        family_hardcopyiii: vl_notype;
        family_hardcopyii: vl_notype;
        family_arriaiigz: vl_notype;
        family_arriaiigx: vl_notype;
        family_stratixiii: vl_notype;
        family_cycloneiii: vl_notype;
        family_cyclone  : vl_notype;
        family_base_cycloneii: vl_notype;
        family_cycloneii: vl_notype;
        family_base_stratix: vl_notype;
        family_base_stratixii: vl_notype;
        family_has_lutram: vl_notype;
        family_has_stratixv_style_ram: vl_notype;
        family_has_stratixiii_style_ram: vl_notype;
        family_has_m512 : vl_notype;
        family_has_megaram: vl_notype;
        family_has_stratixi_style_ram: vl_notype;
        is_write_on_positive_edge: vl_notype;
        lutram_single_port_fast_read: vl_notype;
        lutram_dual_port_fast_read: vl_notype;
        s3_address_aclr_a: vl_notype;
        s3_address_aclr_b: vl_notype;
        i_address_aclr_family_a: vl_notype;
        i_address_aclr_family_b: vl_notype
    );
    port(
        wren_a          : in     vl_logic;
        wren_b          : in     vl_logic;
        rden_a          : in     vl_logic;
        rden_b          : in     vl_logic;
        data_a          : in     vl_logic_vector;
        data_b          : in     vl_logic_vector;
        address_a       : in     vl_logic_vector;
        address_b       : in     vl_logic_vector;
        clock0          : in     vl_logic;
        clock1          : in     vl_logic;
        clocken0        : in     vl_logic;
        clocken1        : in     vl_logic;
        clocken2        : in     vl_logic;
        clocken3        : in     vl_logic;
        aclr0           : in     vl_logic;
        aclr1           : in     vl_logic;
        byteena_a       : in     vl_logic_vector;
        byteena_b       : in     vl_logic_vector;
        addressstall_a  : in     vl_logic;
        addressstall_b  : in     vl_logic;
        q_a             : out    vl_logic_vector;
        q_b             : out    vl_logic_vector;
        eccstatus       : out    vl_logic_vector
    );
    attribute mti_svvh_generic_type : integer;
    attribute mti_svvh_generic_type of width_a : constant is 1;
    attribute mti_svvh_generic_type of widthad_a : constant is 1;
    attribute mti_svvh_generic_type of numwords_a : constant is 1;
    attribute mti_svvh_generic_type of outdata_reg_a : constant is 1;
    attribute mti_svvh_generic_type of address_aclr_a : constant is 1;
    attribute mti_svvh_generic_type of outdata_aclr_a : constant is 1;
    attribute mti_svvh_generic_type of indata_aclr_a : constant is 1;
    attribute mti_svvh_generic_type of wrcontrol_aclr_a : constant is 1;
    attribute mti_svvh_generic_type of byteena_aclr_a : constant is 1;
    attribute mti_svvh_generic_type of width_byteena_a : constant is 1;
    attribute mti_svvh_generic_type of width_b : constant is 1;
    attribute mti_svvh_generic_type of widthad_b : constant is 1;
    attribute mti_svvh_generic_type of numwords_b : constant is 1;
    attribute mti_svvh_generic_type of rdcontrol_reg_b : constant is 1;
    attribute mti_svvh_generic_type of address_reg_b : constant is 1;
    attribute mti_svvh_generic_type of outdata_reg_b : constant is 1;
    attribute mti_svvh_generic_type of outdata_aclr_b : constant is 1;
    attribute mti_svvh_generic_type of rdcontrol_aclr_b : constant is 1;
    attribute mti_svvh_generic_type of indata_reg_b : constant is 1;
    attribute mti_svvh_generic_type of wrcontrol_wraddress_reg_b : constant is 1;
    attribute mti_svvh_generic_type of byteena_reg_b : constant is 1;
    attribute mti_svvh_generic_type of indata_aclr_b : constant is 1;
    attribute mti_svvh_generic_type of wrcontrol_aclr_b : constant is 1;
    attribute mti_svvh_generic_type of address_aclr_b : constant is 1;
    attribute mti_svvh_generic_type of byteena_aclr_b : constant is 1;
    attribute mti_svvh_generic_type of width_byteena_b : constant is 1;
    attribute mti_svvh_generic_type of clock_enable_input_a : constant is 1;
    attribute mti_svvh_generic_type of clock_enable_output_a : constant is 1;
    attribute mti_svvh_generic_type of clock_enable_input_b : constant is 1;
    attribute mti_svvh_generic_type of clock_enable_output_b : constant is 1;
    attribute mti_svvh_generic_type of clock_enable_core_a : constant is 1;
    attribute mti_svvh_generic_type of clock_enable_core_b : constant is 1;
    attribute mti_svvh_generic_type of read_during_write_mode_port_a : constant is 1;
    attribute mti_svvh_generic_type of read_during_write_mode_port_b : constant is 1;
    attribute mti_svvh_generic_type of enable_ecc : constant is 1;
    attribute mti_svvh_generic_type of width_eccstatus : constant is 1;
    attribute mti_svvh_generic_type of ecc_pipeline_stage_enabled : constant is 1;
    attribute mti_svvh_generic_type of operation_mode : constant is 1;
    attribute mti_svvh_generic_type of byte_size : constant is 1;
    attribute mti_svvh_generic_type of read_during_write_mode_mixed_ports : constant is 1;
    attribute mti_svvh_generic_type of ram_block_type : constant is 1;
    attribute mti_svvh_generic_type of init_file : constant is 1;
    attribute mti_svvh_generic_type of init_file_layout : constant is 1;
    attribute mti_svvh_generic_type of maximum_depth : constant is 1;
    attribute mti_svvh_generic_type of intended_device_family : constant is 1;
    attribute mti_svvh_generic_type of lpm_hint : constant is 1;
    attribute mti_svvh_generic_type of lpm_type : constant is 1;
    attribute mti_svvh_generic_type of implement_in_les : constant is 1;
    attribute mti_svvh_generic_type of power_up_uninitialized : constant is 1;
    attribute mti_svvh_generic_type of sim_show_memory_data_in_port_b_layout : constant is 1;
    attribute mti_svvh_generic_type of is_lutram : constant is 3;
    attribute mti_svvh_generic_type of is_bidir_and_wrcontrol_addb_clk0 : constant is 3;
    attribute mti_svvh_generic_type of is_bidir_and_wrcontrol_addb_clk1 : constant is 3;
    attribute mti_svvh_generic_type of check_simultaneous_read_write : constant is 3;
    attribute mti_svvh_generic_type of dual_port_addreg_b_clk0 : constant is 3;
    attribute mti_svvh_generic_type of dual_port_addreg_b_clk1 : constant is 3;
    attribute mti_svvh_generic_type of i_byte_size_tmp : constant is 3;
    attribute mti_svvh_generic_type of i_lutram_read : constant is 3;
    attribute mti_svvh_generic_type of enable_mem_data_b_reading : constant is 3;
    attribute mti_svvh_generic_type of family_arriav : constant is 3;
    attribute mti_svvh_generic_type of family_cyclonev : constant is 3;
    attribute mti_svvh_generic_type of family_base_arriav : constant is 3;
    attribute mti_svvh_generic_type of family_stratixvi : constant is 3;
    attribute mti_svvh_generic_type of family_arriavi : constant is 3;
    attribute mti_svvh_generic_type of family_nightfury : constant is 3;
    attribute mti_svvh_generic_type of family_arriavgz : constant is 3;
    attribute mti_svvh_generic_type of family_stratixv : constant is 3;
    attribute mti_svvh_generic_type of family_hardcopyiv : constant is 3;
    attribute mti_svvh_generic_type of family_hardcopyiii : constant is 3;
    attribute mti_svvh_generic_type of family_hardcopyii : constant is 3;
    attribute mti_svvh_generic_type of family_arriaiigz : constant is 3;
    attribute mti_svvh_generic_type of family_arriaiigx : constant is 3;
    attribute mti_svvh_generic_type of family_stratixiii : constant is 3;
    attribute mti_svvh_generic_type of family_cycloneiii : constant is 3;
    attribute mti_svvh_generic_type of family_cyclone : constant is 3;
    attribute mti_svvh_generic_type of family_base_cycloneii : constant is 3;
    attribute mti_svvh_generic_type of family_cycloneii : constant is 3;
    attribute mti_svvh_generic_type of family_base_stratix : constant is 3;
    attribute mti_svvh_generic_type of family_base_stratixii : constant is 3;
    attribute mti_svvh_generic_type of family_has_lutram : constant is 3;
    attribute mti_svvh_generic_type of family_has_stratixv_style_ram : constant is 3;
    attribute mti_svvh_generic_type of family_has_stratixiii_style_ram : constant is 3;
    attribute mti_svvh_generic_type of family_has_m512 : constant is 3;
    attribute mti_svvh_generic_type of family_has_megaram : constant is 3;
    attribute mti_svvh_generic_type of family_has_stratixi_style_ram : constant is 3;
    attribute mti_svvh_generic_type of is_write_on_positive_edge : constant is 3;
    attribute mti_svvh_generic_type of lutram_single_port_fast_read : constant is 3;
    attribute mti_svvh_generic_type of lutram_dual_port_fast_read : constant is 3;
    attribute mti_svvh_generic_type of s3_address_aclr_a : constant is 3;
    attribute mti_svvh_generic_type of s3_address_aclr_b : constant is 3;
    attribute mti_svvh_generic_type of i_address_aclr_family_a : constant is 3;
    attribute mti_svvh_generic_type of i_address_aclr_family_b : constant is 3;
end altsyncram;

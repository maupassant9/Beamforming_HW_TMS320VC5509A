library verilog;
use verilog.vl_types.all;
entity CYCLONE_PRIM_DFFEAS_HIGH is
    -- This module cannot be connected to from
    -- VHDL because it has unnamed ports.
end CYCLONE_PRIM_DFFEAS_HIGH;
